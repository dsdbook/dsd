module hello;
initial $hello;
endmodule
