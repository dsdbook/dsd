`timescale 1ns/100ps
module name;
reg clk;
reg \clk ;
initial begin
#10 $stop;
end
endmodule
