`timescale 1ns/10ps
module sub(A,B);
input A;
output B;
assign B = A;
endmodule
